module P_Srivastava ();

endmodule