module P_Qian ();

endmodule